`timescale 1ns/1ns

module Controller (input Clk,Start,Rst,Run, input[1:0] stack_out, input is_deque_empty, is_full_X, is_full_Y, is_empty_X, is_empty_Y, is_wall, Finish,
                    output logic our_reset, push, pop_back, pop_front, ld_X, ld_Y, iz_X, iz_Y, sel_X, sel_Y, sel_add, sel_sub, pX_nX, pY_nY, Rd, Wr,
                    output logic Fail, Done, Din, output logic[1:0] dir);




    
endmodule

