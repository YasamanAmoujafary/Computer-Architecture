module Controller(clk, rst, opcode, is_zero,PCWrite, AdrSrc, MemWrite, ResultSrc, ALUControl, ALUSrcA, ALUSrcB,S);
endmodule